
module Global(
 );
reg [31:0] reg_array [31:0];

endmodule